module Not(
    input in,
    output out
);

    assign out = ~in;
endmodule
module Not(
    input in,
    output out
);

    assign out = ~a;
endmodule